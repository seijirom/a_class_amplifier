* Z:\HOME\ANAGIX\WORK\YSS_PMOS\A_CLASS_AMPLIFIER\AMP_HARUNA.ASC
M13 N010 N009 N004 N001 PMOS L=10U W=27000U
R3 N001 N009 10K
R4 N009 0 20K
R5 N002 N004 30
R6 N001 N002 3K
R7 N010 0 4.5K
M14 0 N010 N005 N001 PMOS L=10U W=1800U
R8 N001 N005 10K
M15 N006 N003 N001 N001 PMOS L=10U W=45000U
M16 N003 N003 N001 N001 PMOS L=10U W=1800U
R13 N003 0 1K
M17 0 N005 N006 N001 PMOS L=10U W=45000U
*C1 N001 N002 {100U}
*C2 N009 N008 {100U}
*C3 N007 N006 {1000U}
*V1 N001 0 10
*V2 N008 0 SINE 0 0.11 1K AC 1
*R1 N007 0 8
.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\ANAGIX\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
* .STEP PARAM R1K LIST  100K 200K
*.INCLUDE MODELS/PMOS
* 2020/08/18 VER1.1 CGS0 CGD0 CJ
* BSIM3 MODEL 
* BY C.TAKAHASHI

.MODEL YSS_PMOS PMOS
+ LEVEL = 49
+ VERSION = 3.3
+ PARAMCHK = 1
+ BINUNIT = 1
+ MOBMOD = 1
+ CAPMOD = 3
+ NOIMOD = 1
+ VTH0 = _0.9
+ K1 = 0.53
+ K2 = _0.0186
+ K3 = 80
+ K3B = 0
+ W0 = 4.5E_06
+ NLX = 1.74E_007
+ VBM = _3
+ DVT0 = 5.2
+ DVT1 = 0.53
+ DVT2 = _0.032
+ DVT0W = 0
+ DVT1W = 5300000
+ DVT2W = _0.032
+ U0 = 600
+ UA = 2.25E_9
+ UB = 5.87E_19
+ UC = 0 
+ VSAT = 90000
+ A0 = 0.00
+ AGS = 0.0
+ B0 = 0
+ B1 = 0
+ KETA = _0.047
+ A1 = 1
+ A2 = 0
+ RDSW = 30K 
+ PRWG = 0
+ PRWB = 0
+ WR = 1
+ LINT = 1.3E_6
+ WINT = 0
+ DWG = 0
+ DWB = 0
+ VOFF = _0.5
+ NFACTOR = 0
+ ETA0 = 0.08
+ ETAB = _0.07
+ DSUB = 0.56
+ CIT = 0
+ CDSC = 0.00024
+ CDSCD = 0
+ CDSCB = 0
+ PCLM = 10
+ PDIBLC1 = 0
+ PDIBLC2 = 0.02
+ PDIBLCB = 0
+ DROUT = 0.56
+ PVAG = 0
#+ PSCBE1 = 0
+ PSCBE2 = 2E_4
+ DELTA = 0.01
+ NGATE = 0
+ ALPHA0 = 0
+ ALPHA1 = 0
+ BETA0 = 30
+ RSH = 0
+ XPART = 0
+ CGSO = 1.22E_9
+ CGDO = 1.22E_9
+ CJ   = 2.04E_8
+ MJ   = 0.5
+ CJSWG = 5E_010
+ MJSWG = 0.33
+ PBSWG = 1
+ CGSL = 0
+ CGDL = 0
+ CKAPPA = 0.6
+ CLC = 1E_007
+ CLE = 0.6
+ DLC = 0
+ DWC = 0
+ WL = 0
+ WLN = 1
+ WW = 0
+ WWN = 1
+ WWL = 0
+ LL = 0
+ LLN = 1
+ LW = 0
+ LWN = 1
+ LWL = 0
+ TNOM = 27
+ UTE = _1.5
+ KT1 = _0.11
+ KT1L = 0
+ KT2 = _0.022
+ UA1 = 4.31E_009
+ UB1 = _7.61E_018
+ UC1 = _5.6E_011
+ AT = 33000
+ PRT = 0
+ NOIA = 9.9E+18
+ NOIB = 2.4E3
+ NOIC = 1.4E_012
+ EM = 41000000
+ AF = 1
+ EF = 1
+ KF = 0
+ TOX = 6E_08
+ XJ = 1.5E_007
+ NCH = 1.7E+017
+ NSUB = 6E+016
+ XT = 1.55E_007
+ BINUNIT = 1
.TRAN 10M
.STEP PARAM L20 10U 60U 10U
.BACKANNO
.END
